// $Id: $
// File name:   fifobuff.sv
// Created:     3/24/2015
// Author:      Andy Shi
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: fifo for operations

module fifobuff(
input wire clk, n_rst, read_date,
input reg [2:0] opcode_in,
output reg [2:0] opcode_out
);

endmodule