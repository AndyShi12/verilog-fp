// $Id: $
// File name:   wrapper.sv
// Created:     4/22/2015
// Author:      Kyunghoon Jung
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Wrapper file for floating point co-processor
