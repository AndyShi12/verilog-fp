// $Id: $
// File name:   tb_addsub.sv
// Created:     3/28/2015
// Author:      Andy Shi
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: test bench for add/sub
`timescale 1ns/10ps

module tb_addsub();

localparam	CLK_PERIOD	= 2.5;
localparam	CHECK_DELAY = 1; 
